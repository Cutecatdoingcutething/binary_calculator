library ieee ;
use ieee.std_logic_1164.ALL ;
use ieee.std_logic_arith.ALL ;
use ieee.std_logic_unsigned.ALL ;

package state_package is
	type state_type is (S1, S2, S3, S4, S5, S6, S7) ;
end package ;

package body state_package is
end package body ;